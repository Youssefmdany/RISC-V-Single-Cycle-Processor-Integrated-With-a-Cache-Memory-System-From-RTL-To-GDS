

parameter R_Type   = 7'b0110011;
parameter I_Type_1 = 7'b0000011;
parameter I_Type_2 = 7'b0010011;
parameter I_Type_3 = 7'b1100111;
parameter S_Type   = 7'b0100011;
parameter U_Type_1 = 7'b0010111;
parameter U_Type_2 = 7'b0110111;
parameter J_Type   = 7'b1101111;
parameter B_Type   = 7'b1100011;



